module FPGA_CLOCK_tb;
        AX_DEBOUNCE_tb ax_debounce_tb_ ();
        BEEP_tb beep_tb_ ();
        SEG_tb seg_tb_ ();
        SQUARE_WAVE_GENERATOR_tb sw_gen_tb_ ();
        TIME_MODULE_tb_1 time_module_tb_ ();
        TIME_MODULE_tb_2 time_module_tb__ ();
        TIME_SEG_UNIT_tb time_seg_unit_tb_ ();
        TIMER_tb timer_tb_ ();
endmodule
